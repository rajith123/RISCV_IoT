`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module ALU(
  input         clock,
  input         reset,
  input  [3:0]  io_fn,
  input  [31:0] io_in2,
  input  [31:0] io_in1,
  output [31:0] io_out,
  output [31:0] io_adder_out
);
  wire  _T_12;
  wire [32:0] _T_14;
  wire [32:0] _T_15;
  wire [31:0] _T_16;
  wire [31:0] _T_17;
  wire [32:0] _T_18;
  wire [31:0] sum;
  wire  _T_19;
  wire  _T_20;
  wire  _T_21;
  wire  _T_22;
  wire  _T_23;
  wire  _T_26;
  wire  less;
  wire [4:0] shamt;
  wire  _T_27;
  wire  _T_28;
  wire  _T_29;
  wire [15:0] _T_34;
  wire [31:0] _T_35;
  wire [15:0] _T_36;
  wire [31:0] _GEN_0;
  wire [31:0] _T_37;
  wire [31:0] _T_39;
  wire [31:0] _T_40;
  wire [23:0] _T_44;
  wire [31:0] _GEN_1;
  wire [31:0] _T_45;
  wire [23:0] _T_46;
  wire [31:0] _GEN_2;
  wire [31:0] _T_47;
  wire [31:0] _T_49;
  wire [31:0] _T_50;
  wire [27:0] _T_54;
  wire [31:0] _GEN_3;
  wire [31:0] _T_55;
  wire [27:0] _T_56;
  wire [31:0] _GEN_4;
  wire [31:0] _T_57;
  wire [31:0] _T_59;
  wire [31:0] _T_60;
  wire [29:0] _T_64;
  wire [31:0] _GEN_5;
  wire [31:0] _T_65;
  wire [29:0] _T_66;
  wire [31:0] _GEN_6;
  wire [31:0] _T_67;
  wire [31:0] _T_69;
  wire [31:0] _T_70;
  wire [30:0] _T_74;
  wire [31:0] _GEN_7;
  wire [31:0] _T_75;
  wire [30:0] _T_76;
  wire [31:0] _GEN_8;
  wire [31:0] _T_77;
  wire [31:0] _T_79;
  wire [31:0] _T_80;
  wire [31:0] shin;
  wire  _T_82;
  wire  _T_83;
  wire [32:0] _T_84;
  wire [32:0] _T_85;
  wire [32:0] _T_86;
  wire [31:0] shout_r;
  wire [15:0] _T_91;
  wire [31:0] _T_92;
  wire [15:0] _T_93;
  wire [31:0] _GEN_9;
  wire [31:0] _T_94;
  wire [31:0] _T_96;
  wire [31:0] _T_97;
  wire [23:0] _T_101;
  wire [31:0] _GEN_10;
  wire [31:0] _T_102;
  wire [23:0] _T_103;
  wire [31:0] _GEN_11;
  wire [31:0] _T_104;
  wire [31:0] _T_106;
  wire [31:0] _T_107;
  wire [27:0] _T_111;
  wire [31:0] _GEN_12;
  wire [31:0] _T_112;
  wire [27:0] _T_113;
  wire [31:0] _GEN_13;
  wire [31:0] _T_114;
  wire [31:0] _T_116;
  wire [31:0] _T_117;
  wire [29:0] _T_121;
  wire [31:0] _GEN_14;
  wire [31:0] _T_122;
  wire [29:0] _T_123;
  wire [31:0] _GEN_15;
  wire [31:0] _T_124;
  wire [31:0] _T_126;
  wire [31:0] _T_127;
  wire [30:0] _T_131;
  wire [31:0] _GEN_16;
  wire [31:0] _T_132;
  wire [30:0] _T_133;
  wire [31:0] _GEN_17;
  wire [31:0] _T_134;
  wire [31:0] _T_136;
  wire [31:0] shout_l;
  wire  _T_137;
  wire [31:0] _T_138;
  wire  _T_139;
  wire [31:0] _T_140;
  wire  _T_141;
  wire [31:0] _T_142;
  wire [31:0] _T_143;
  wire [31:0] _T_144;
  wire [31:0] bitwise_logic;
  wire  _T_145;
  wire  _T_146;
  wire  _T_147;
  wire  _T_148;
  wire  _T_149;
  wire  _T_150;
  wire  _T_154;
  wire [31:0] _T_155;
  wire [31:0] _T_156;
  wire [31:0] _T_157;
  wire [31:0] out_xpr_length;
  assign io_out = out_xpr_length;
  assign io_adder_out = sum;
  assign _T_12 = io_fn[3];
  assign _T_14 = 32'h0 - io_in2;
  assign _T_15 = $unsigned(_T_14);
  assign _T_16 = _T_15[31:0];
  assign _T_17 = _T_12 ? _T_16 : io_in2;
  assign _T_18 = io_in1 + _T_17;
  assign sum = _T_18[31:0];
  assign _T_19 = io_in1[31];
  assign _T_20 = io_in2[31];
  assign _T_21 = _T_19 == _T_20;
  assign _T_22 = sum[31];
  assign _T_23 = io_fn[0];
  assign _T_26 = _T_23 ? _T_20 : _T_19;
  assign less = _T_21 ? _T_22 : _T_26;
  assign shamt = io_in2[4:0];
  assign _T_27 = io_fn == 4'h5;
  assign _T_28 = io_fn == 4'hd;
  assign _T_29 = _T_27 | _T_28;
  assign _T_34 = io_in1[31:16];
  assign _T_35 = {{16'd0}, _T_34};
  assign _T_36 = io_in1[15:0];
  assign _GEN_0 = {{16'd0}, _T_36};
  assign _T_37 = _GEN_0 << 16;
  assign _T_39 = _T_37 & 32'hffff0000;
  assign _T_40 = _T_35 | _T_39;
  assign _T_44 = _T_40[31:8];
  assign _GEN_1 = {{8'd0}, _T_44};
  assign _T_45 = _GEN_1 & 32'hff00ff;
  assign _T_46 = _T_40[23:0];
  assign _GEN_2 = {{8'd0}, _T_46};
  assign _T_47 = _GEN_2 << 8;
  assign _T_49 = _T_47 & 32'hff00ff00;
  assign _T_50 = _T_45 | _T_49;
  assign _T_54 = _T_50[31:4];
  assign _GEN_3 = {{4'd0}, _T_54};
  assign _T_55 = _GEN_3 & 32'hf0f0f0f;
  assign _T_56 = _T_50[27:0];
  assign _GEN_4 = {{4'd0}, _T_56};
  assign _T_57 = _GEN_4 << 4;
  assign _T_59 = _T_57 & 32'hf0f0f0f0;
  assign _T_60 = _T_55 | _T_59;
  assign _T_64 = _T_60[31:2];
  assign _GEN_5 = {{2'd0}, _T_64};
  assign _T_65 = _GEN_5 & 32'h33333333;
  assign _T_66 = _T_60[29:0];
  assign _GEN_6 = {{2'd0}, _T_66};
  assign _T_67 = _GEN_6 << 2;
  assign _T_69 = _T_67 & 32'hcccccccc;
  assign _T_70 = _T_65 | _T_69;
  assign _T_74 = _T_70[31:1];
  assign _GEN_7 = {{1'd0}, _T_74};
  assign _T_75 = _GEN_7 & 32'h55555555;
  assign _T_76 = _T_70[30:0];
  assign _GEN_8 = {{1'd0}, _T_76};
  assign _T_77 = _GEN_8 << 1;
  assign _T_79 = _T_77 & 32'haaaaaaaa;
  assign _T_80 = _T_75 | _T_79;
  assign shin = _T_29 ? io_in1 : _T_80;
  assign _T_82 = shin[31];
  assign _T_83 = _T_12 & _T_82;
  assign _T_84 = {_T_83,shin};
  assign _T_85 = $signed(_T_84);
  assign _T_86 = $signed(_T_85) >>> shamt;
  assign shout_r = _T_86[31:0];
  assign _T_91 = shout_r[31:16];
  assign _T_92 = {{16'd0}, _T_91};
  assign _T_93 = shout_r[15:0];
  assign _GEN_9 = {{16'd0}, _T_93};
  assign _T_94 = _GEN_9 << 16;
  assign _T_96 = _T_94 & 32'hffff0000;
  assign _T_97 = _T_92 | _T_96;
  assign _T_101 = _T_97[31:8];
  assign _GEN_10 = {{8'd0}, _T_101};
  assign _T_102 = _GEN_10 & 32'hff00ff;
  assign _T_103 = _T_97[23:0];
  assign _GEN_11 = {{8'd0}, _T_103};
  assign _T_104 = _GEN_11 << 8;
  assign _T_106 = _T_104 & 32'hff00ff00;
  assign _T_107 = _T_102 | _T_106;
  assign _T_111 = _T_107[31:4];
  assign _GEN_12 = {{4'd0}, _T_111};
  assign _T_112 = _GEN_12 & 32'hf0f0f0f;
  assign _T_113 = _T_107[27:0];
  assign _GEN_13 = {{4'd0}, _T_113};
  assign _T_114 = _GEN_13 << 4;
  assign _T_116 = _T_114 & 32'hf0f0f0f0;
  assign _T_117 = _T_112 | _T_116;
  assign _T_121 = _T_117[31:2];
  assign _GEN_14 = {{2'd0}, _T_121};
  assign _T_122 = _GEN_14 & 32'h33333333;
  assign _T_123 = _T_117[29:0];
  assign _GEN_15 = {{2'd0}, _T_123};
  assign _T_124 = _GEN_15 << 2;
  assign _T_126 = _T_124 & 32'hcccccccc;
  assign _T_127 = _T_122 | _T_126;
  assign _T_131 = _T_127[31:1];
  assign _GEN_16 = {{1'd0}, _T_131};
  assign _T_132 = _GEN_16 & 32'h55555555;
  assign _T_133 = _T_127[30:0];
  assign _GEN_17 = {{1'd0}, _T_133};
  assign _T_134 = _GEN_17 << 1;
  assign _T_136 = _T_134 & 32'haaaaaaaa;
  assign shout_l = _T_132 | _T_136;
  assign _T_137 = io_fn == 4'h7;
  assign _T_138 = io_in1 & io_in2;
  assign _T_139 = io_fn == 4'h6;
  assign _T_140 = io_in1 | io_in2;
  assign _T_141 = io_fn == 4'h4;
  assign _T_142 = io_in1 ^ io_in2;
  assign _T_143 = _T_141 ? _T_142 : io_in1;
  assign _T_144 = _T_139 ? _T_140 : _T_143;
  assign bitwise_logic = _T_137 ? _T_138 : _T_144;
  assign _T_145 = io_fn == 4'h0;
  assign _T_146 = io_fn == 4'h8;
  assign _T_147 = _T_145 | _T_146;
  assign _T_148 = io_fn == 4'ha;
  assign _T_149 = io_fn == 4'hb;
  assign _T_150 = _T_148 | _T_149;
  assign _T_154 = io_fn == 4'h1;
  assign _T_155 = _T_154 ? shout_l : bitwise_logic;
  assign _T_156 = _T_29 ? shout_r : _T_155;
  assign _T_157 = _T_150 ? {{31'd0}, less} : _T_156;
  assign out_xpr_length = _T_147 ? sum : _T_157;
endmodule
